// class env_configs extens uvm_object;
//     `uvm_object_utils(env_configs)

   

// endclass